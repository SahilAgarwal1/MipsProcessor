library ieee;
use ieee.std_logic_1164.all;

package gen_mux_package is
    type mux_array is array (natural range <>) of std_logic_vector(31 downto 0);
end package;

package body gen_mux_package is
end package body;
